module d_ff(clk,q,rst,d); 
input d,clk,rst; 
output reg q; 
always@(posedge clk) 
begin 
if(rst==1) 
q=1'b0;  
else 
q=d; 
end 
endmodule
